`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/07/2022 08:42:44 PM
// Design Name: 
// Module Name: sevdectwelvehr
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sevdectwelvehr(a_in,out);
  input [7:0] a_in;
  output reg [13:0] out;
    always @(*) begin
        case (a_in)
            8'b00000000: out = 14'b00000010000001;//00
            8'b00000001: out = 14'b00000011001111;//01
            8'b00000010: out = 14'b00000010010010;//02
            8'b00000011: out = 14'b00000010000110;//03
            8'b00000100: out = 14'b00000011001100;//04
            8'b00000101: out = 14'b00000010100100;//05
            8'b00000110: out = 14'b00000010100000;//06
            8'b00000111: out = 14'b00000010001111;//07
            8'b00001000: out = 14'b00000010000000;//08
            8'b00001001: out = 14'b00000010000100;//09
            8'b00010000: out = 14'b10011110000001;//10
            8'b00010001: out = 14'b10011111001111;//11
            8'b00010010: out = 14'b10011110010010;//12
            8'b00010011: out = 14'b00000011001111;//01
            8'b00010100: out = 14'b00000010010010;//02
            8'b00010101: out = 14'b00000010000110;//03
            8'b00010110: out = 14'b00000011001100;//04
            8'b00010111: out = 14'b00000010100100;//05
            8'b00011000: out = 14'b00000010100000;//06
            8'b00011001: out = 14'b00000010001111;//07
            8'b00100000: out = 14'b00000010000000;//08
            8'b00100001: out = 14'b00000010000100;//09
            8'b00100010: out = 14'b10011110000001;//10
            8'b00100011: out = 14'b10011111001111;//11
            8'b00100100: out = 14'b00000010000001;//00
         endcase
       end           
endmodule


